//------------------------------------------------------------------------------
//File       : dummy_dut.sv
//Author     : Nirvara Reddy/1BM23EC170
//Created    : 2026-02-10
//Module     : dummy_dut
//Project    : SystemVerilog and Verification (23EC6PE2SV)
//Faculty    : Prof. Ajaykumar Devarapalli
//Description: A placeholder dummy DUT for the class-based Packet verification lab.
//------------------------------------------------------------------------------

module dummy_dut;
endmodule
